LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.ALL;

ENTITY Decode IS
    PORT (
        clk : IN STD_LOGIC;
        reset : IN STD_LOGIC;
        MemRead_EXCUTESTAGE : IN STD_LOGIC;
        RD_EXCUTESTAGE : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
        InputPC : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        Instruction : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        INPORTDATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
        RFData1,RFData2 : IN std_logic_vector(31 DOWNTO 0);
        RD1, RD2, ImmValue : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
        RS1, RS2, RD : OUT STD_LOGIC_VECTOR(2 DOWNTO 0);
        ControlSignals : OUT STD_LOGIC_VECTOR(24 DOWNTO 0);
        HazardSignal : OUT STD_LOGIC);
END ENTITY Decode;

ARCHITECTURE Decode OF Decode IS
    COMPONENT ControlUnit IS
        PORT (
            clk, reset : IN STD_LOGIC;
            opCode : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
            SignalVector : OUT STD_LOGIC_VECTOR(24 DOWNTO 0));
    END COMPONENT ControlUnit;

    COMPONENT mux2 IS
        GENERIC (n : INTEGER := 1);
        PORT (
            IN1, IN2 : IN STD_LOGIC_VECTOR(n - 1 DOWNTO 0);
            SEl : IN STD_LOGIC;
            OUT1 : OUT STD_LOGIC_VECTOR(n - 1 DOWNTO 0));
    END COMPONENT mux2;

    COMPONENT HazardDU IS
        PORT (
            clk : IN STD_LOGIC;
            MemRead : IN STD_LOGIC;
            RS1, RS2, RD : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
            hazard1 : OUT STD_LOGIC);
    END COMPONENT HazardDU;
    SIGNAL OpCode : STD_LOGIC_VECTOR(5 DOWNTO 0);
    SIGNAL Reg1Add : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL Reg2Add : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL Reg1Data : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL Reg2Data : STD_LOGIC_VECTOR(31 DOWNTO 0);
    SIGNAL CONTSIG : STD_LOGIC_VECTOR(24 DOWNTO 0);

    -----------------------------------------------------------------------------------------
    --CONTROL UNIT SIGNALS-------------------------
    SIGNAL RegWrite : STD_LOGIC := '0';
    SIGNAL InPort : STD_LOGIC := '0';
    SIGNAL OutPort : STD_LOGIC := '0';
    SIGNAL RegImm : STD_LOGIC := '0';
    SIGNAL RegDst : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    SIGNAL ALUOp : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
    SIGNAL JmpCond : STD_LOGIC_VECTOR(1 DOWNTO 0) := "00";
    SIGNAL Branch : STD_LOGIC := '0';
    SIGNAL SpHeap : STD_LOGIC := '0';
    SIGNAL MemWrite : STD_LOGIC := '0';
    SIGNAL MemRead : STD_LOGIC := '0';
    SIGNAL MemAluToReg : STD_LOGIC := '0';
    SIGNAL PcRd2 : STD_LOGIC := '0';
    SIGNAL PcMem : STD_LOGIC := '0';
    SIGNAL HLT : STD_LOGIC := '0';
    SIGNAL SWAP : STD_LOGIC := '0';
    SIGNAL SWInt : STD_LOGIC := '0';
    SIGNAL RTISIg : STD_LOGIC := '0';
    SIGNAL Flush : STD_LOGIC := '0';
    SIGNAL HWINT : STD_LOGIC := '0';
    --HAZARD SIGNAL----------------------------
    SIGNAL hazardSig : STD_LOGIC := '0';

BEGIN

    CU : ControlUnit PORT MAP(clk => clk, reset => reset, opCode => Opcode, signalVector => CONTSIG);
    -- INPORTREG: my_nDFF GENERIC MAP(32) PORT MAP(clk=>clk,Rst=>reset,en=>'0',d=>(OTHERS=>'0'),q=>INPORTDATA);
    INPORTMUX : mux2 GENERIC MAP(32) PORT MAP(SEl => InPort, IN1 => RFData1, IN2 => INPORTDATA, OUT1 => RD1);
    HDU : HazardDU PORT MAP(clk => clk, MemRead => MemRead_EXCUTESTAGE, RS1 => Reg1Add, RS2 => Reg2Add, RD => RD_EXCUTESTAGE, hazard1 => hazardSig);
    HDUMUX : mux2 GENERIC MAP(25) PORT MAP(SEl => hazardSig, IN1 => CONTSIG, IN2 => (OTHERS => '0'), OUT1 => ControlSignals);
    InPort <= CONTSIG(22);
    Opcode <= Instruction(31 DOWNTO 26);
    Reg1Add <= Instruction(25 DOWNTO 23);
    Reg2Add <= Instruction(22 DOWNTO 20);
    ImmValue <= x"0000" & Instruction(15 DOWNTO 0);
    RS1 <= Instruction(25 DOWNTO 23);
    RS2 <= Instruction(22 DOWNTO 20);
    RD <= Instruction(19 DOWNTO 17);
    RD2 <=RFData2;
    HazardSignal <= hazardSig;

END Decode;