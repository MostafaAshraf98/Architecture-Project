LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY Integration IS
    PORT ();
END ENTITY;
ARCHITECTURE a_Integration OF Integration IS
BEGIN

END ARCHITECTURE;