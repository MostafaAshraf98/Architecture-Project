LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY Execute_Unit IS
    PORT ();
END ENTITY;
ARCHITECTURE a_Execute_Unit OF Execute_Unit IS
BEGIN

END ARCHITECTURE;